`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/11/13 21:02:21
// Design Name: 
// Module Name: instruction
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instruction(addr, instruction);
	input [31:0] addr;
	output [31:0] instruction;
	reg [31:0] instruction;
	reg [31:0] InsMem[0:63];
	integer i;
	initial begin
		InsMem[0]  = 32'b00100000000010000000000000100000; //addi $t0, $zero, 0x20
		InsMem[1]  = 32'b00100000000010010000000000100111; //addi $t1, $zero, 0x27
		InsMem[2]  = 32'b00000001000010011000000000100100; //and $s0, $t0, $t1
		InsMem[3]  = 32'b00000001000010011000000000100101; //or $s0, $t0, $t1
		InsMem[4]  = 32'b10101100000100000000000000000100; //sw $s0, 4($zero)
		InsMem[5]  = 32'b10101100000010000000000000001000; //sw $t0, 8($zero)
		InsMem[6]  = 32'b00000001000010011000100000100000; //add $s1, $t0, $t1
		InsMem[7]  = 32'b00000001000010011001000000100010; //sub $s2, $t0, $t1
		InsMem[8]  = 32'b00010010001100100000000000001001; //beq $s1, $s2, error0
		InsMem[9]  = 32'b10001100000100010000000000000100; //lw $s1, 4($zero)
		InsMem[10] = 32'b00110010001100100000000000011000; //andi $s2, $s1, 0x18
		InsMem[11] = 32'b00010010001100100000000000001001; //beq $s1, $s2, error1
		InsMem[12] = 32'b10001100000100110000000000001000; //lw $s3, 8($zero)
		InsMem[13] = 32'b00010010000100110000000000001010; //beq $s0, $s3, error2
		InsMem[14] = 32'b00000010010100011010000000101010; //slt $s4, $s2, $s1 (Last)
		InsMem[15] = 32'b00010010100000000000000000001111; //beq $s4, $0, EXIT
		InsMem[16] = 32'b00000010001000001001000000100000; //add $s2, $s1, $0
		InsMem[17] = 32'b00001000000000000000000000001110; //j Last
		InsMem[18] = 32'b00100000000010000000000000000000; //addi $t0, $0, 0(error0)
		InsMem[19] = 32'b00100000000010010000000000000000; //addi $t1, $0, 0
		InsMem[20] = 32'b00001000000000000000000000011111; //j EXIT
		InsMem[21] = 32'b00100000000010000000000000000001; //addi $t0, $0, 1(error1)
		InsMem[22] = 32'b00100000000010010000000000000001; //addi $t1, $0, 1
		InsMem[23] = 32'b00001000000000000000000000011111; //j EXIT
		InsMem[24] = 32'b00100000000010000000000000000010; //addi $t0, $0, 2(error2)
		InsMem[25] = 32'b00100000000010010000000000000010; //addi $t1, $0, 2
		InsMem[26] = 32'b00001000000000000000000000011111; //j EXIT
		InsMem[27] = 32'b00100000000010000000000000000011; //addi $t0, $0, 3(error3)
		InsMem[28] = 32'b00100000000010010000000000000011; //addi $t1, $0, 3
		InsMem[29] = 32'b00001000000000000000000000011111; //j EXIT
	end
	
	always @ (addr)
	begin
		instruction = InsMem[addr[7:0]>>2];
	end
endmodule


